LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY Execute IS
	PORT( Read_data1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			Read_data2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ALU_Result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END Execute;

ARCHITECTURE behavior OF Execute IS

BEGIN
	ALU_Result <= read_data1 + read_data2;
END behavior;